module controlUnit  (
    input wire [5:0]  instr_op , 
    output wire reg_dst      ,   
    output wire  branch    ,     
    output wire  mem_read ,  
    output wire  mem_to_reg  ,
    output wire [1:0]  alu_op  ,        
    output wire  mem_write  , 
    output wire  alu_src     ,    
    output wire  reg_write  , 
    );

// ------------------------------
// Insert your solution below
// ------------------------------ 

endmodule
